-----------------------------------------------------------------------------
--
--  Conway TB constants package
--
--  This package defines constant vectors used in the conway test bench
--
--  Revision History
--     03/15/2019 Sundar Pandian       Initial version
--
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

use work.constants.all;

package TBConstants is

	constant NumTests : integer := 5; -- number of tests

	-- test vector array
    type TestVector is array(NumTests-1 downto 0, ARRYSIZE*ARRYSIZE-1 downto 0) of std_logic;

    constant InputTest : TestVector := (

	   ('0', '0', '0', '0', '0', '0', '1', '0', '0', '0', 
		'1', '0', '0', '0', '0', '1', '0', '0', '1', '0', 
		'0', '0', '0', '1', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '1', '0', '0', '0', '1', '0', '1', 
		'1', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '1', '0', '1', '0', '1', '0', '0', 
		'0', '0', '0', '0', '0', '1', '0', '0', '0', '0', 
		'0', '1', '0', '0', '0', '0', '0', '0', '1', '1'),

	   ('0', '1', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '1', '0', '0', '1', '0', '1', '0', 
		'0', '1', '0', '1', '0', '0', '0', '0', '1', '0', 
		'1', '0', '1', '0', '1', '0', '0', '0', '1', '0', 
		'0', '0', '0', '1', '1', '0', '0', '0', '1', '0', 
		'0', '0', '1', '0', '0', '0', '0', '0', '0', '1', 
		'0', '0', '1', '0', '0', '0', '0', '1', '1', '0', 
		'1', '0', '0', '0', '0', '0', '1', '1', '0', '0', 
		'1', '0', '0', '0', '0', '1', '0', '0', '1', '1', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0'),

	   ('0', '0', '1', '0', '0', '1', '0', '1', '0', '1', 
		'0', '1', '0', '0', '0', '1', '1', '0', '1', '0', 
		'0', '0', '0', '0', '0', '1', '0', '0', '0', '0', 
		'0', '0', '0', '1', '0', '0', '0', '0', '0', '1', 
		'0', '0', '0', '0', '0', '0', '0', '1', '0', '1', 
		'0', '0', '1', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '1', '0', '1', '0', '0', '0', '0', '0', 
		'0', '0', '1', '0', '0', '0', '1', '0', '1', '0', 
		'0', '0', '0', '1', '0', '0', '0', '0', '0', '0', 
		'1', '0', '0', '1', '0', '0', '1', '0', '1', '0'),

	   ('0', '0', '0', '0', '0', '1', '0', '0', '0', '1', 
		'0', '0', '1', '0', '0', '0', '0', '0', '1', '0', 
		'0', '0', '0', '0', '0', '0', '1', '0', '0', '0', 
		'0', '0', '0', '0', '1', '0', '0', '1', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '1', '0', '0', '0', '0', '0', '0', '1', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '1', '1', '1', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'1', '0', '0', '0', '1', '0', '0', '0', '0', '1'),

	   ('0', '0', '0', '0', '1', '0', '0', '0', '0', '1', 
		'1', '0', '0', '0', '1', '0', '0', '1', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'1', '0', '0', '0', '0', '0', '0', '0', '1', '0', 
		'0', '0', '0', '0', '0', '1', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '1', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '1', '1', '0', 
		'0', '0', '0', '0', '0', '0', '0', '1', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '1', '0', 
		'0', '1', '0', '0', '0', '1', '0', '0', '0', '1')
    );

    constant OutputTest : TestVector := (

	   ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0'),

	   ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '1', '0', '0', '0', '0', '0', 
		'0', '0', '0', '1', '1', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '1', '0', '0', '1', '0', '1', '1', '0', 
		'0', '1', '0', '1', '0', '1', '1', '1', '1', '1', 
		'0', '0', '1', '1', '0', '0', '0', '0', '0', '1', 
		'0', '0', '0', '0', '1', '1', '1', '0', '1', '1', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0'),

	   ('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '1', '1', '1', '1', '1', 
		'0', '0', '0', '0', '0', '1', '1', '1', '1', '0', 
		'0', '0', '1', '0', '0', '0', '1', '0', '0', '0', 
		'0', '1', '0', '1', '0', '0', '0', '0', '0', '0', 
		'1', '1', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0'),

	   ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0'),

	   ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '1', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '1', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '1', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0')
    );

end package TBConstants;